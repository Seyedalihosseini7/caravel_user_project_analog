magic
tech sky130A
timestamp 1633983915
<< nwell >>
rect -9000 0 -6000 3000
<< pdiff >>
rect -8900 2860 -6100 2900
rect -8900 1740 -8860 2860
rect -6140 1740 -6100 2860
rect -8900 1700 -6100 1740
rect -8900 1260 -6100 1300
rect -8900 140 -8860 1260
rect -6140 140 -6100 1260
rect -8900 100 -6100 140
<< pdiffc >>
rect -8860 1740 -6140 2860
rect -8860 140 -6140 1260
<< nsubdiff >>
rect -8900 1580 -6100 1600
rect -8900 1420 -8880 1580
rect -6120 1420 -6100 1580
rect -8900 1400 -6100 1420
<< nsubdiffcont >>
rect -8880 1420 -6120 1580
<< locali >>
rect -9000 2860 -6000 2900
rect -9000 1740 -8860 2860
rect -6140 1740 -6000 2860
rect -9000 1700 -6000 1740
rect -9000 1580 -6000 1600
rect -9000 1420 -8880 1580
rect -6120 1420 -6000 1580
rect -9000 1400 -6000 1420
rect -9000 1260 -6000 1300
rect -9000 140 -8860 1260
rect -6140 140 -6000 1260
rect -9000 100 -6000 140
<< viali >>
rect -6300 1850 -6250 2750
rect -8850 1450 -8750 1550
rect -6300 250 -6250 1150
<< metal1 >>
rect -8900 1550 -8700 3000
rect -8900 1450 -8850 1550
rect -8750 1450 -8700 1550
rect -8900 0 -8700 1450
rect -6400 2750 -6200 3000
rect -6400 1850 -6300 2750
rect -6250 1850 -6200 2750
rect -6400 1150 -6200 1850
rect -6400 250 -6300 1150
rect -6250 250 -6200 1150
rect -6400 0 -6200 250
<< end >>
